----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:08:50 12/01/2016 
-- Design Name: 
-- Module Name:    DataMem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DataMem is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (31 downto 0);
           din : in  STD_LOGIC_VECTOR (31 downto 0);
           dout : out  STD_LOGIC_VECTOR (31 downto 0);
           selwr : in  STD_LOGIC;		
           selrd : in  STD_LOGIC);
			  
--			  m8: out std_logic_vector(31 downto 0);
--			  m9: out std_logic_vector(31 downto 0);
--			  m10: out std_logic_vector(31 downto 0);
--			  m11: out std_logic_vector(31 downto 0);
--			  m12: out std_logic_vector(31 downto 0));		
end DataMem;

architecture Behavioral of DataMem is
TYPE ram IS ARRAY (0 TO 35) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
signal mem : ram := ram'(x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000",x"00000000",x"00000000");

signal mem1 : ram := ram'(x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
								x"00000000",x"00000000",x"00000000");
								
signal memaddr : std_logic_vector(31 downto 0);

begin

--process(clk, rst, selrd, selwr, addr)
--begin
----if(clk'event and clk = '0') then
--if (rst = '0') then
--	if (selrd = '1' or selwr = '1') then
--		memaddr <= addr;
--	else
--		memaddr <= x"00000000";
--	end if;
--end if;
----end if;
--end process;

process(clk, rst, selwr, addr, din)
begin
if(clk'event and clk = '0') then
	if(rst = '0') then
		if(selwr = '1') then
			mem(conv_integer(addr)) <= din;
		end if;
	else
		mem <= mem1;
	end if;
end if;	
end process;

process(rst, selrd, addr, mem)
begin
if (clk = '0') then
	if (rst = '0') then
		if (selrd = '1') then
			dout <= mem(conv_integer(addr));
		--else
			dout <= x"00000000";
		end if;
		--dout <= x"00000000";
	end if;
--	dout <= x"00000000";
end if;
end process;

--m8<=mem(8);
--m9<=mem(9);
--m10<=mem(10);
--m11<=mem(11);
--m12<=mem(12);
							
--TYPE ram IS ARRAY (0 TO 35) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
--signal s_arr_temp : ram := ram'("10110111111000010101000101100011", "01010110000110001001011000111000", "11110100010100000100010011010101",
--"10010010100001111011111010001110", "00110000101111110011100001000111", "11001110111101101011001000000000",
--"01101101001011100010101110111001", "00001011011001011010010101110010", "10101001100111010001111100101011",
--"01000111110101001001100011100100", "11100110000011000001001010011101", "10000100010000111000110001010110",
--"00100010011110110000011000001111", "11000000101100100111111111001000", "01011110111010011111100110000001",
--"11111101001000010111001100111010", "10011011010110001110110011110011", "00111001100100000110011010101100",
--"11010111110001111110000001100101", "01110101111111110101101000011110", "00010100001101101101001111010111",
--"10110010011011100100110110010000", "01010000101001011100011101001001", "11101110110111010100000100000010",
--"10001101000101001011101010111011", "00101011010011000011010001110100", "00000000000000000000000000000000",
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000",
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000",
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000");
----signal din : STD_LOGIC_VECTOR (31 downto 0);
--signal s_arr_temp1 : ram := ram'("10110111111000010101000101100011", "01010110000110001001011000111000", "11110100010100000100010011010101",
--"10010010100001111011111010001110", "00110000101111110011100001000111", "11001110111101101011001000000000",
--"01101101001011100010101110111001", "00001011011001011010010101110010", "10101001100111010001111100101011",
--"01000111110101001001100011100100", "11100110000011000001001010011101", "10000100010000111000110001010110",
--"00100010011110110000011000001111", "11000000101100100111111111001000", "01011110111010011111100110000001",
--"11111101001000010111001100111010", "10011011010110001110110011110011", "00111001100100000110011010101100",
--"11010111110001111110000001100101", "01110101111111110101101000011110", "00010100001101101101001111010111",
--"10110010011011100100110110010000", "01010000101001011100011101001001", "11101110110111010100000100000010",
--"10001101000101001011101010111011", "00101011010011000011010001110100", "00000000000000000000000000000000",
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000",
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000",
--"00000000000000000000000000000000", "00000000000000000000000000000000", "00000000000000000000000000000000");
--
--
--begin
--
--process(clk, rst, addr, selwr, selrd, din)
--begin
--  if(clk'event and clk = '1') then
--	 if(rst = '0') then
--		if(selwr = '1') then
--		s_arr_temp(conv_integer(addr)) <= din;
--		elsif(selrd = '1') then
--		dout <= s_arr_temp(conv_integer(addr));
--		end if;
--	else--if(rst = '1') then
--	s_arr_temp <= s_arr_temp1;
--	end if;
--  end if;
--end process;




end Behavioral;